`timescale 1ns/1ps  

module APB_Slave (
    // glob
    input logic PCLK,
    input logic PRESET,

    // APB Inferface Signals
    input logic [3:0] PADDR,
    input logic PWRITE,
    input logic PSEL,
    input logic PENABLE,
    input logic [31:0] PWDATA,
    output logic [31:0] PRDATA,
    output logic PREADY
);

    logic [31:0] slv_reg0, slv_reg1, slv_reg2, slv_reg3;

    always_ff @( posedge PCLK, posedge PRESET ) begin
        if (PRESET) begin
            slv_reg0 <= 32'b0;
            slv_reg1 <= 32'b0;
            slv_reg2 <= 32'b0;
            slv_reg3 <= 32'b0;
        end else begin
            PREADY <= 1'b0;
            if (PSEL && PENABLE) begin
                // w/o wait states
                PREADY <= 1'b1;
                if (PWRITE) begin
                    case (PADDR[3:2])
                        2'd0: slv_reg0 <= PWDATA;
                        2'd1: slv_reg1 <= PWDATA;
                        2'd2: slv_reg2 <= PWDATA;
                        2'd3: slv_reg3 <= PWDATA;
                    endcase
                end else begin
                    case (PADDR[3:2])
                        2'd0: PRDATA <= slv_reg0;
                        2'd1: PRDATA <= slv_reg1;
                        2'd2: PRDATA <= slv_reg2;
                        2'd3: PRDATA <= slv_reg3;
                    endcase
                end
            end
        end
    end
endmodule
