`timescale 1ns / 1ps

module APB_GPO (
    // global signals
    input  logic        PCLK,
    input  logic        PRESET,
    // APB Interface Signals
    input  logic [ 2:0] PADDR,
    input  logic        PWRITE,
    input  logic        PSEL,
    input  logic        PENABLE,
    input  logic [31:0] PWDATA,
    output logic [31:0] PRDATA,
    output logic        PREADY,
    // external signals ports
    output logic [ 3:0] gpo
);

    logic [3:0] mode;
    logic [3:0] out_data;

    APB_Slave_GPO_Interface U_APB_GPO_Intf (.*);
    apb_gpo U_GPO (.*);

endmodule


module APB_Slave_GPO_Interface (
    // global signals
    input  logic        PCLK,
    input  logic        PRESET,
    // APB Interface Signals
    input  logic [ 2:0] PADDR,
    input  logic        PWRITE,
    input  logic        PSEL,
    input  logic        PENABLE,
    input  logic [31:0] PWDATA,
    output logic [31:0] PRDATA,
    output logic        PREADY,
    // internal signals
    output logic [ 3:0] mode,
    output logic [ 3:0] out_data
);
    logic [31:0] slv_reg0, slv_reg1;  //, slv_reg2, slv_reg3;

    assign mode = slv_reg0[3:0];
    assign out_data = slv_reg1[3:0];

    always_ff @(posedge PCLK, posedge PRESET) begin
        if (PRESET) begin
            slv_reg0 <= 0;
            slv_reg1 <= 0;
            // slv_reg2 <= 0;
            // slv_reg3 <= 0;
        end else begin
            PREADY <= 1'b0;
            if (PSEL & PENABLE) begin
                PREADY <= 1'b1;
                if (PWRITE) begin
                    case (PADDR[2]) 
                        1'd0: slv_reg0 <= PWDATA;   // 0x00
                        1'd1: slv_reg1 <= PWDATA;   // 0x04
                        // 2'd2: slv_reg2 <= PWDATA;
                        // 2'd3: slv_reg3 <= PWDATA;
                    endcase
                end else begin
                    case (PADDR[2])
                        1'd0: PRDATA <= slv_reg0;
                        1'd1: PRDATA <= slv_reg1;
                        // 2'd2: PRDATA <= slv_reg2;
                        // 2'd3: PRDATA <= slv_reg3;
                    endcase

                end
            end
        end
    end
endmodule

// mode: 1 - output enabled, 0 - high impedance
module apb_gpo (
    input  logic [3:0] mode,
    input  logic [3:0] out_data,
    output logic [3:0] gpo
);

    genvar i;

    generate
        for (i = 0; i < 4; i++) begin
            assign gpo[i] = mode[i] ? out_data[i] : 1'bz;
        end
    endgenerate

endmodule
